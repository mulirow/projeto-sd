module rx(clk1, in, ledData, recorder);
    input clk1, in;
    output [7:0]ledData;
    output reg [3:0]recorder;

    

endmodule
